module emblem_gen(
    input wire [9:0] x,
    input wire [9:0] y,
    input wire active,
    output reg draw,
    output reg [5:0] rgb
);

    localparam [9:0] EMBLEM_X0 = 240;
    localparam [9:0] EMBLEM_X1 = 400;
    localparam [9:0] EMBLEM_Y0 = 144;
    localparam [9:0] EMBLEM_Y1 = 320;
    localparam [9:0] EMBLEM_CENTER_X = (EMBLEM_X0 + EMBLEM_X1) >> 1;

    localparam [5:0] COLOR_BLACK = 6'b000000;
    localparam [5:0] COLOR_GOLD = 6'b110110;
    localparam [5:0] COLOR_RED = 6'b100100;
    localparam [5:0] COLOR_WHITE = 6'b111111;

    localparam [9:0] BORDER_THICKNESS = 3;
    localparam [9:0] CHEVRON_BORDER_THICK = 3;

    // Chevron parameters
    // Original bitmap: 85 pixels wide, 100 pixels tall
    // Scaled 2x for display: 170 pixels wide, 200 pixels tall
    localparam [9:0] CHEVRON_BITMAP_WIDTH = 85;
    localparam [9:0] CHEVRON_BITMAP_HEIGHT = 100;
    localparam [9:0] CHEVRON_SCALE = 2;  // 2x scale
    localparam [9:0] CHEVRON_WIDTH = CHEVRON_BITMAP_WIDTH * CHEVRON_SCALE;  // 170 pixels
    localparam [9:0] CHEVRON_HEIGHT = CHEVRON_BITMAP_HEIGHT * CHEVRON_SCALE;  // 200 pixels
    localparam [9:0] CHEVRON_X = EMBLEM_CENTER_X - (CHEVRON_WIDTH >> 1);
    localparam [9:0] CHEVRON_Y = EMBLEM_Y0 - 14;  // Positioned at top of emblem, moved up 4 pixels
    localparam [6:0] CHEVRON_BITMAP_MIN_ROW = 7'd37;
    localparam [6:0] CHEVRON_BITMAP_MAX_ROW = 7'd76;

    localparam integer LION_WIDTH_PIX = 48;
    localparam [9:0] LION_WIDTH = 48;
    localparam [9:0] LION_HEIGHT = 45;
    localparam [9:0] TOP_LION_Y = EMBLEM_Y0 + 16;
    localparam [9:0] BOTTOM_LION_Y = EMBLEM_Y0 + 112;
    localparam [9:0] LEFT_LION_X = EMBLEM_X0 + 18;  // Moved 2 pixels left to increase spacing
    localparam [9:0] RIGHT_LION_X = EMBLEM_X1 - 18 - LION_WIDTH;  // Moved 2 pixels right to increase spacing
    localparam [9:0] CENTER_LION_X = EMBLEM_CENTER_X - (LION_WIDTH >> 1);

    function automatic [LION_WIDTH_PIX-1:0] lion_row;
        input [5:0] idx;
        begin
            case (idx)
                6'd0:  lion_row = 48'h00001C000000;
                6'd1:  lion_row = 48'h00001FC00000;
                6'd2:  lion_row = 48'h2000FFE00000;
                6'd3:  lion_row = 48'h3202FFF00000;
                6'd4:  lion_row = 48'h3A01FFFC00E0;
                6'd5:  lion_row = 48'h3F81FFFCC1F8;
                6'd6:  lion_row = 48'h3FC7FFF8C1FC;
                6'd7:  lion_row = 48'h1FE1FF99C1F8;
                6'd8:  lion_row = 48'h1FF1FFFFC3FC;
                6'd9:  lion_row = 48'h0FF3FFC007FE;
                6'd10: lion_row = 48'h01F7FFF01FF0;
                6'd11: lion_row = 48'h30F1FFCCBFF8;
                6'd12: lion_row = 48'h3071FFFFFF90;
                6'd13: lion_row = 48'h3F33FFFFFF80;
                6'd14: lion_row = 48'h3F33FFFFFF80;
                6'd15: lion_row = 48'h1FE07FFFFF00;
                6'd16: lion_row = 48'h0FE07FFFFD00;
                6'd17: lion_row = 48'h03C0FFFFF800;
                6'd18: lion_row = 48'h31801FFFFC00;
                6'd19: lion_row = 48'h39803FFFFC00;
                6'd20: lion_row = 48'h3F003FFFFE00;
                6'd21: lion_row = 48'h1F002FFFEF80;
                6'd22: lion_row = 48'h0E003FC07FFC;
                6'd23: lion_row = 48'h0E00FFFFFFFE;
                6'd24: lion_row = 48'h0C01FFFFFFFC;
                6'd25: lion_row = 48'h0C07FFFFFFFF;
                6'd26: lion_row = 48'h080FFFFA4FFF;
                6'd27: lion_row = 48'h081FFE0088FC;
                6'd28: lion_row = 48'h0C3FFF8000F8;
                6'd29: lion_row = 48'h0C3FFFF80058;
                6'd30: lion_row = 48'h071FFFFE0000;
                6'd31: lion_row = 48'h03FFFFFE0000;
                6'd32: lion_row = 48'h003FFFFF0000;
                6'd33: lion_row = 48'h0007FEFF0000;
                6'd34: lion_row = 48'h0007FEFF0000;
                6'd35: lion_row = 48'h0007FEFF0000;
                6'd36: lion_row = 48'h007FFE7F0000;
                6'd37: lion_row = 48'h00FFFC7F8C00;
                6'd38: lion_row = 48'h01FFE07FDE00;
                6'd39: lion_row = 48'h01FF403FFE00;
                6'd40: lion_row = 48'h01FF001BFF00;
                6'd41: lion_row = 48'h01FF0009FF80;
                6'd42: lion_row = 48'h00FF00007E00;
                6'd43: lion_row = 48'h003F8C007E00;
                6'd44: lion_row = 48'h0017FC006200;
                default: lion_row = 48'h000000000000;
            endcase
        end
    endfunction

    wire is_lion_pixel;
    reg [5:0] lion_col_offset;
    reg [5:0] lion_row_offset;
    reg lion_box_hit;

    always @(*) begin
        reg [9:0] temp_col;
        reg [9:0] temp_row;
        
        lion_box_hit = 0;
        lion_col_offset = 0;
        lion_row_offset = 0;
        temp_col = 0;
        temp_row = 0;

        // Check if the pixel is within the Y-range of the top two lions
        if (y >= TOP_LION_Y && y < (TOP_LION_Y + LION_HEIGHT)) begin
            // Check for top-left lion
            if (x >= LEFT_LION_X && x < (LEFT_LION_X + LION_WIDTH)) begin
                temp_col = x - LEFT_LION_X;
                temp_row = y - TOP_LION_Y;
                lion_col_offset = temp_col[5:0];
                lion_row_offset = temp_row[5:0];
                lion_box_hit = 1;
            // Check for top-right lion
            end else if (x >= RIGHT_LION_X && x < (RIGHT_LION_X + LION_WIDTH)) begin
                temp_col = x - RIGHT_LION_X;
                temp_row = y - TOP_LION_Y;
                lion_col_offset = temp_col[5:0];
                lion_row_offset = temp_row[5:0];
                lion_box_hit = 1;
            end
        // Check if the pixel is within the Y-range of the bottom lion
        end else if (y >= BOTTOM_LION_Y && y < (BOTTOM_LION_Y + LION_HEIGHT)) begin
            // Check for bottom lion
            if (x >= CENTER_LION_X && x < (CENTER_LION_X + LION_WIDTH)) begin
                temp_col = x - CENTER_LION_X;
                temp_row = y - BOTTOM_LION_Y;
                lion_col_offset = temp_col[5:0];
                lion_row_offset = temp_row[5:0];
                lion_box_hit = 1;
            end
        end
    end

    // Look up the pixel from the bitmap ROM only if it was inside one of the lion boxes
    wire [LION_WIDTH_PIX-1:0] lion_mask;
    assign lion_mask = lion_row(lion_row_offset[5:0]);
    assign is_lion_pixel = lion_box_hit ? lion_mask[lion_col_offset[5:0]] : 1'b0;

    // Rows are stored relative to CHEVRON_BITMAP_MIN_ROW to drop the zero padding above/below the chevron.
    function automatic [95:0] chevron_row;
        input [5:0] idx;
        begin
            case (idx)
                6'd0:  chevron_row = 96'h000000000020000000000000;  // row 37
                6'd1:  chevron_row = 96'h000000000070000000000000;  // row 38
                6'd2:  chevron_row = 96'h0000000000F8000000000000;  // row 39
                6'd3:  chevron_row = 96'h0000000001FC000000000000;  // row 40
                6'd4:  chevron_row = 96'h0000000003FE000000000000;  // row 41
                6'd5:  chevron_row = 96'h0000000007FF000000000000;  // row 42
                6'd6:  chevron_row = 96'h000000000FFF800000000000;  // row 43
                6'd7:  chevron_row = 96'h000000001FFFC00000000000;  // row 44
                6'd8:  chevron_row = 96'h000000003FFFE00000000000;  // row 45
                6'd9:  chevron_row = 96'h000000007FFFF00000000000;  // row 46
                6'd10: chevron_row = 96'h00000000FFDFF80000000000;  // row 47
                6'd11: chevron_row = 96'h00000001FF8FFC0000000000;  // row 48
                6'd12: chevron_row = 96'h00000003FF07FE0000000000;  // row 49
                6'd13: chevron_row = 96'h00000007FE03FF0000000000;  // row 50
                6'd14: chevron_row = 96'h0000000FFC01FF8000000000;  // row 51
                6'd15: chevron_row = 96'h0000001FF800FFC000000000;  // row 52
                6'd16: chevron_row = 96'h0000003FF0007FE000000000;  // row 53
                6'd17: chevron_row = 96'h0000007FE0003FF000000000;  // row 54
                6'd18: chevron_row = 96'h000000FFC0001FF800000000;  // row 55
                6'd19: chevron_row = 96'h000001FF80000FFC00000000;  // row 56
                6'd20: chevron_row = 96'h000003FF000007FE00000000;  // row 57
                6'd21: chevron_row = 96'h000007FE000003FF00000000;  // row 58
                6'd22: chevron_row = 96'h00000FFC000001FF80000000;  // row 59
                6'd23: chevron_row = 96'h00001FF8000000FFC0000000;  // row 60
                6'd24: chevron_row = 96'h00003FF00000007FE0000000;  // row 61
                6'd25: chevron_row = 96'h00007FE00000003FF0000000;  // row 62
                6'd26: chevron_row = 96'h0000FFC00000001FF8000000;  // row 63
                6'd27: chevron_row = 96'h0001FF800000000FFC000000;  // row 64
                6'd28: chevron_row = 96'h0003FF0000000007FE000000;  // row 65
                6'd29: chevron_row = 96'h0007FE0000000003FF000000;  // row 66
                6'd30: chevron_row = 96'h000FFC0000000001FF800000;  // row 67
                6'd31: chevron_row = 96'h001FF80000000000FFC00000;  // row 68
                6'd32: chevron_row = 96'h003FF000000000007FE00000;  // row 69
                6'd33: chevron_row = 96'h001FE000000000003FC00000;  // row 70
                6'd34: chevron_row = 96'h000FC000000000001F800000;  // row 71
                6'd35: chevron_row = 96'h000F8000000000000F800000;  // row 72
                6'd36: chevron_row = 96'h000F00000000000007800000;  // row 73
                6'd37: chevron_row = 96'h000E00000000000003800000;  // row 74
                6'd38: chevron_row = 96'h000C00000000000001800000;  // row 75
                6'd39: chevron_row = 96'h000800000000000000800000;  // row 76
                default: chevron_row = 96'h000000000000000000000000;
            endcase
        end
    endfunction

    wire is_chevron_pixel;
    reg [6:0] chevron_scaled_col;
    reg [6:0] chevron_scaled_row;
    reg chevron_box_hit;
    wire chevron_row_in_range;

    always @(*) begin
        reg [9:0] temp_scaled_col;
        reg [9:0] temp_scaled_row;
        
        chevron_box_hit = 1'b0;
        chevron_scaled_col = 0;
        chevron_scaled_row = 0;
        temp_scaled_col = 0;
        temp_scaled_row = 0;

        // Check if the pixel is within the chevron bounds (scaled)
        if (y >= CHEVRON_Y && y < (CHEVRON_Y + CHEVRON_HEIGHT) &&
            x >= CHEVRON_X && x < (CHEVRON_X + CHEVRON_WIDTH)) begin
            // Scale down to original bitmap coordinates (divide by scale factor)
            temp_scaled_col = (x - CHEVRON_X) >> 1;
            temp_scaled_row = (y - CHEVRON_Y) >> 1;
            chevron_scaled_col = temp_scaled_col[6:0];
            chevron_scaled_row = temp_scaled_row[6:0];
            chevron_box_hit = 1;
        end
    end

    wire [6:0] chevron_row_idx;
    wire [6:0] chevron_bit_idx;
    wire [95:0] chevron_mask;
    
    assign chevron_row_in_range = (chevron_scaled_row >= CHEVRON_BITMAP_MIN_ROW) && (chevron_scaled_row <= CHEVRON_BITMAP_MAX_ROW);
    assign chevron_row_idx = chevron_scaled_row - CHEVRON_BITMAP_MIN_ROW;
    assign chevron_bit_idx = 7'd95 - chevron_scaled_col[6:0];
    assign chevron_mask = chevron_row_in_range ? chevron_row(chevron_row_idx[5:0]) : 96'h0;
    assign is_chevron_pixel = (chevron_box_hit && chevron_row_in_range) ? chevron_mask[chevron_bit_idx] : 1'b0;

    // Chevron border detection: check if pixel is within 3 pixels of a chevron pixel
    // Helper function to check if a pixel at (px, py) is a chevron pixel
    function automatic is_chevron_at;
        input [9:0] px;
        input [9:0] py;
        reg [9:0] p_col_offset, p_row_offset;
        reg [6:0] p_scaled_col, p_scaled_row;
        reg p_box_hit;
        reg p_row_in_range;
        reg [6:0] p_row_idx, p_bit_idx;
        reg [95:0] p_mask;
        begin
            is_chevron_at = 1'b0;
            if (py >= CHEVRON_Y && py < (CHEVRON_Y + CHEVRON_HEIGHT) &&
                px >= CHEVRON_X && px < (CHEVRON_X + CHEVRON_WIDTH)) begin
                p_col_offset = (px - CHEVRON_X) >> 1;
                p_row_offset = (py - CHEVRON_Y) >> 1;
                p_scaled_col = p_col_offset[6:0];
                p_scaled_row = p_row_offset[6:0];
                p_row_in_range = (p_scaled_row >= CHEVRON_BITMAP_MIN_ROW) && 
                                 (p_scaled_row <= CHEVRON_BITMAP_MAX_ROW);
                p_row_idx = p_scaled_row - CHEVRON_BITMAP_MIN_ROW;
                p_bit_idx = 7'd95 - p_scaled_col[6:0];
                p_mask = p_row_in_range ? chevron_row(p_row_idx[5:0]) : 96'h0;
                is_chevron_at = p_row_in_range ? p_mask[p_bit_idx] : 1'b0;
            end
        end
    endfunction

    // Check all pixels within Manhattan distance 3 (7x7 grid = 49 pixels, but only check those within distance 3)
    reg is_chevron_border;
    reg border_found;
    
    always @(*) begin
        reg nearby_is_chevron;
        
        border_found = 1'b0;
        is_chevron_border = 1'b0;
        nearby_is_chevron = 1'b0;
        
        // Only check for border if we're in the expanded chevron region and not a chevron pixel
        if (!is_chevron_pixel &&
            y >= (CHEVRON_Y > CHEVRON_BORDER_THICK ? CHEVRON_Y - CHEVRON_BORDER_THICK : 0) && 
            y < (CHEVRON_Y + CHEVRON_HEIGHT + CHEVRON_BORDER_THICK) &&
            x >= (CHEVRON_X > CHEVRON_BORDER_THICK ? CHEVRON_X - CHEVRON_BORDER_THICK : 0) && 
            x < (CHEVRON_X + CHEVRON_WIDTH + CHEVRON_BORDER_THICK)) begin
            
            // Check all offsets within Manhattan distance 3
            // dx=-3: dy can be 0
            if (x >= 3 && !border_found) begin
                nearby_is_chevron = is_chevron_at(x - 3, y);
                if (nearby_is_chevron) border_found = 1'b1;
            end
            
            // dx=-2: dy can be 0, 1
            if (!border_found && x >= 2) begin
                nearby_is_chevron = is_chevron_at(x - 2, y) || is_chevron_at(x - 2, y - 1) || 
                                    is_chevron_at(x - 2, y + 1);
                if (nearby_is_chevron) border_found = 1'b1;
            end
            
            // dx=-1: dy can be 0, 1, 2
            if (!border_found && x >= 1) begin
                nearby_is_chevron = is_chevron_at(x - 1, y) || is_chevron_at(x - 1, y - 1) || 
                                    is_chevron_at(x - 1, y + 1) || is_chevron_at(x - 1, y - 2) || 
                                    is_chevron_at(x - 1, y + 2);
                if (nearby_is_chevron) border_found = 1'b1;
            end
            
            // dx=0: dy can be 1, 2, 3
            if (!border_found) begin
                nearby_is_chevron = is_chevron_at(x, y - 1) || is_chevron_at(x, y + 1) || 
                                    is_chevron_at(x, y - 2) || is_chevron_at(x, y + 2) ||
                                    is_chevron_at(x, y - 3) || is_chevron_at(x, y + 3);
                if (nearby_is_chevron) border_found = 1'b1;
            end
            
            // dx=+1: dy can be 0, 1, 2
            if (!border_found) begin
                nearby_is_chevron = is_chevron_at(x + 1, y) || is_chevron_at(x + 1, y - 1) || 
                                    is_chevron_at(x + 1, y + 1) || is_chevron_at(x + 1, y - 2) || 
                                    is_chevron_at(x + 1, y + 2);
                if (nearby_is_chevron) border_found = 1'b1;
            end
            
            // dx=+2: dy can be 0, 1
            if (!border_found) begin
                nearby_is_chevron = is_chevron_at(x + 2, y) || is_chevron_at(x + 2, y - 1) || 
                                    is_chevron_at(x + 2, y + 1);
                if (nearby_is_chevron) border_found = 1'b1;
            end
            
            // dx=+3: dy can be 0
            if (!border_found) begin
                nearby_is_chevron = is_chevron_at(x + 3, y);
                if (nearby_is_chevron) border_found = 1'b1;
            end
        end
        
        is_chevron_border = border_found;
    end

    function automatic [6:0] shield_width;
        input [7:0] y_addr;
        begin
            shield_width = 7'd78;

            if (y_addr < 8'd88) begin
                shield_width = (y_addr < 8'd83) ? 7'd77 : 7'd76;
            end else if (y_addr < 8'd96) begin
                shield_width = (y_addr < 8'd92) ? 7'd75 : 7'd74;
            end else if (y_addr < 8'd99) begin
                shield_width = 7'd73;
            end else if (y_addr < 8'd102) begin
                shield_width = 7'd72;
            end else if (y_addr < 8'd105) begin
                shield_width = 7'd71;
            end else if (y_addr < 8'd108) begin
                shield_width = 7'd70;
            end else if (y_addr < 8'd111) begin
                shield_width = 7'd69;
            end else if (y_addr < 8'd114) begin
                shield_width = 7'd68;
            end else if (y_addr < 8'd117) begin
                shield_width = 7'd67;
            end else if (y_addr < 8'd120) begin
                shield_width = 7'd66;
            end else if (y_addr < 8'd123) begin
                shield_width = 7'd65;
            end else if (y_addr < 8'd126) begin
                shield_width = 7'd64;
            end else if (y_addr < 8'd128) begin
                shield_width = 7'd63;
            end else if (y_addr < 8'd130) begin
                shield_width = 7'd62;
            end else if (y_addr < 8'd132) begin
                shield_width = 7'd61;
            end else if (y_addr < 8'd134) begin
                shield_width = 7'd60;
            end else if (y_addr < 8'd136) begin
                shield_width = 7'd59;
            end else if (y_addr < 8'd138) begin
                shield_width = 7'd58;
            end else if (y_addr < 8'd140) begin
                shield_width = 7'd57;
            end else if (y_addr < 8'd142) begin
                shield_width = 7'd56;
            end else if (y_addr < 8'd144) begin
                shield_width = 7'd55;
            end else if (y_addr < 8'd146) begin
                shield_width = 7'd54;
            end else if (y_addr < 8'd156) begin
                shield_width = 7'd53 - 7'(y_addr - 8'd146);
            end else begin
                shield_width = 7'd42 - 7'((y_addr - 8'd156) << 1);
            end
        end
    endfunction

    reg draw_flag;

    always @(*) begin
        reg [6:0] half_width;
        reg [6:0] inner_half;
        reg shield_border;
        reg [9:0] abs_dx;
        reg [9:0] rel_y;

        half_width = 0;
        inner_half = 0;
        shield_border = 0;
        draw_flag = 0;
        rgb = 6'b000000;
        abs_dx = (x >= EMBLEM_CENTER_X) ? (x - EMBLEM_CENTER_X) : (EMBLEM_CENTER_X - x);
        rel_y = y - EMBLEM_Y0;

        if (active && (y >= EMBLEM_Y0) && (y < EMBLEM_Y1)) begin
            half_width = shield_width(rel_y[7:0]);
            if (abs_dx <= {3'b0, half_width}) begin
                draw_flag = 1;
                rgb = COLOR_GOLD;

                inner_half = (half_width > BORDER_THICKNESS[6:0]) ? (half_width - BORDER_THICKNESS[6:0]) : 7'b0;
                if ((abs_dx > {3'b0, inner_half}) || (rel_y < BORDER_THICKNESS)) shield_border = 1;

                if (is_chevron_border) rgb = COLOR_BLACK;
                if (is_chevron_pixel) rgb = COLOR_WHITE;
                if (is_lion_pixel) rgb = COLOR_RED;
                if (shield_border) rgb = COLOR_BLACK;
            end
        end
        draw = draw_flag;
    end

endmodule
